library verilog;
use verilog.vl_types.all;
entity tb_mux2x1 is
end tb_mux2x1;
