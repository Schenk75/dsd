library verilog;
use verilog.vl_types.all;
entity testbench_comb is
end testbench_comb;
