library verilog;
use verilog.vl_types.all;
entity tb_Encoder8x3 is
end tb_Encoder8x3;
