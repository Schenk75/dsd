library verilog;
use verilog.vl_types.all;
entity comb_prim is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end comb_prim;
