library verilog;
use verilog.vl_types.all;
entity tb_mux4x1 is
end tb_mux4x1;
