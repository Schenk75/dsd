library verilog;
use verilog.vl_types.all;
entity tb_comb_Y2 is
end tb_comb_Y2;
